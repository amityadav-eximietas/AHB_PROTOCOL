/////////////////////////////////////////////////////////////////
//  file name     : ahb_master_pkg.sv
//  owner name    : amit yadav & anupam mathur
//  module name   : ahb masterter package
//  company name  : eximietas design
//////////////////////////////////////////////////////////////////

`ifndef AHB_MASTER_PKG_SV
`define AHB_MASTER_PKG_SV

`include "ahb_master_if.sv"

package ahb_master_pkg;
   import uvm_pkg::*;
endpackage

`endif //AHB_MASTER_PKG_SV

