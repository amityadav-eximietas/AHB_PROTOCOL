/////////////////////////////////////////////////////////////////
//  file name     : ahb_env_pkg.sv
//  owner name    : amit yadav & anupam mathur
//  module name   : ahb environment package
//  company name  : eximietas design
//////////////////////////////////////////////////////////////////

`ifndef AHB_ENV_PKG_SV
`define AHB_ENV_PKG_SV
`include "ahb_master_if.sv"
`include "ahb_slave_if.sv"

package ahb_env_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
    
  `include "ahb_defines.svh"
  `include "ahb_seq_item.sv"
  
  `include "ahb_master_config.svh" 
  `include "ahb_master_driver.sv"
  `include "ahb_master_seqr.sv"
  `include "ahb_master_monitor.sv"
  `include "ahb_master_agent.sv"
  `include "ahb_master_base_seqs.sv"

  `include "ahb_slave_seq_item.sv"
  `include "ahb_slave_config.svh"
  `include "ahb_common_object.sv"
  `include "ahb_slave_driver.sv"
  `include "ahb_slave_monitor.sv"
  `include "ahb_slave_agent.sv"
  

  `include "ahb_env_config.svh"
  `include "ahb_scoreboard.sv"	
  `include "ahb_env.sv"  
endpackage

`endif //AHB_ENV_PKG_SV

